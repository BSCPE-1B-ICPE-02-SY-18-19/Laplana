CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 10 6 120 10
176 80 1534 813
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 976 37 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5130 0 0
2
5.89883e-315 0
0
2 +V
167 294 256 0 1 3
0 14
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
43529.7 0
0
7 Pulser~
4 93 306 0 10 12
0 18 19 15 20 0 0 5 5 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3124 0 0
2
43529.7 1
0
9 CC 7-Seg~
183 1052 322 0 17 19
10 9 8 7 6 5 4 3 21 2
2 2 2 2 2 2 2 2
0
0 0 21104 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3421 0 0
2
43529.7 2
0
9 2-In AND~
219 684 215 0 3 22
0 16 10 17
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8157 0 0
2
43529.7 3
0
9 2-In AND~
219 438 168 0 3 22
0 13 12 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
43529.7 4
0
6 74112~
219 759 270 0 7 32
0 14 17 15 17 14 22 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8901 0 0
2
43529.7 5
0
6 74112~
219 610 353 0 7 32
0 14 16 15 16 14 10 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
7361 0 0
2
43529.7 6
0
6 74112~
219 431 459 0 7 32
0 14 13 15 13 14 23 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
4747 0 0
2
43529.7 7
0
6 74112~
219 243 551 0 7 32
0 14 14 15 14 14 24 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
972 0 0
2
43529.7 8
0
6 74LS48
188 961 515 0 14 29
0 11 10 12 13 25 26 3 4 5
6 7 8 9 27
0
0 0 4848 0
6 74LS48
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
43529.7 9
0
38
1 9 0 0 0 0 0 1 4 0 0 4
976 45
976 272
1052 272
1052 280
7 7 0 0 0 0 0 11 4 0 0 3
993 479
1067 479
1067 358
8 6 0 0 0 0 0 11 4 0 0 3
993 488
1061 488
1061 358
9 5 0 0 0 0 0 11 4 0 0 3
993 497
1055 497
1055 358
10 4 0 0 0 0 0 11 4 0 0 3
993 506
1049 506
1049 358
11 3 0 0 0 0 0 11 4 0 0 3
993 515
1043 515
1043 358
12 2 0 0 0 0 0 11 4 0 0 3
993 524
1037 524
1037 358
13 1 0 0 0 0 0 11 4 0 0 3
993 533
1031 533
1031 358
6 0 10 0 0 4096 0 8 0 0 11 2
640 335
641 335
0 1 11 0 0 4224 0 0 11 15 0 5
798 299
798 443
894 443
894 479
929 479
0 2 10 0 0 8320 0 0 11 30 0 5
641 297
641 452
902 452
902 488
929 488
0 3 12 0 0 8320 0 0 11 28 0 5
483 300
483 458
908 458
908 497
929 497
0 4 13 0 0 8320 0 0 11 38 0 5
333 300
333 467
915 467
915 506
929 506
0 1 14 0 0 4096 0 0 2 25 0 5
295 300
256 300
256 273
294 273
294 265
7 0 11 0 0 0 0 7 0 0 0 4
783 234
798 234
798 299
811 299
1 0 14 0 0 0 0 2 0 0 20 2
294 265
294 265
0 0 14 0 0 4096 0 0 0 20 23 2
355 265
355 373
1 1 14 0 0 8192 0 8 7 0 0 5
610 290
610 265
729 265
729 207
759 207
1 1 14 0 0 8320 0 9 8 0 0 4
431 396
431 265
610 265
610 290
1 1 14 0 0 4096 0 10 9 0 0 4
243 488
243 265
431 265
431 396
5 5 14 0 0 0 0 8 7 0 0 4
610 365
610 356
759 356
759 282
5 5 14 0 0 16384 0 9 8 0 0 6
431 471
431 489
384 489
384 356
610 356
610 365
5 5 14 0 0 0 0 10 9 0 0 6
243 563
355 563
355 373
476 373
476 471
431 471
3 0 15 0 0 8192 0 3 0 0 35 4
117 297
140 297
140 398
206 398
4 2 14 0 0 12416 0 10 10 0 0 8
219 533
219 578
295 578
295 300
256 300
256 478
219 478
219 515
2 0 16 0 0 4096 0 8 0 0 27 4
586 317
563 317
563 297
548 297
0 4 16 0 0 4224 0 0 8 29 0 3
548 200
548 335
586 335
2 7 12 0 0 0 0 6 9 0 0 5
414 177
414 205
483 205
483 423
455 423
3 1 16 0 0 0 0 6 5 0 0 4
459 168
548 168
548 206
660 206
2 7 10 0 0 0 0 5 8 0 0 6
660 224
652 224
652 297
641 297
641 317
634 317
2 0 17 0 0 8192 0 7 0 0 32 4
735 234
722 234
722 299
712 299
3 4 17 0 0 8320 0 5 7 0 0 6
705 215
712 215
712 299
712 299
712 252
735 252
3 0 15 0 0 0 0 8 0 0 35 3
580 326
554 326
554 399
3 0 15 0 0 0 0 9 0 0 35 3
401 432
397 432
397 399
3 3 15 0 0 20608 0 10 7 0 0 8
213 524
206 524
206 398
242 398
242 399
702 399
702 243
729 243
1 0 13 0 0 0 0 6 0 0 37 3
414 159
367 159
367 300
4 0 13 0 0 0 0 9 0 0 38 3
407 441
367 441
367 300
7 2 13 0 0 0 0 10 9 0 0 6
267 515
333 515
333 300
367 300
367 423
407 423
3
-35 0 0 0 700 0 0 0 0 3 2 1 2
15 Chintzy CPU BRK
0 0 0 51
23 102 964 146
29 109 957 141
51 4 - bit synchronous counter waveform timing diagram
-21 0 0 0 700 0 0 0 0 3 2 1 2
15 Chintzy CPU BRK
0 0 0 9
64 66 199 94
72 72 190 92
9 BSCpE 1-B
-21 0 0 0 700 0 0 0 0 3 2 1 2
15 Chintzy CPU BRK
0 0 0 17
63 47 275 75
72 53 265 73
17 Laplana, Larry C.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
